`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:39:52 04/17/2019 
// Design Name: 
// Module Name:    Structural 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Structural(
    input s1,
    input s0,
    input i0,
    input i1,
    input i2,
    input i3,
    output d
    );


endmodule
